library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

-- author: CZW
-- date: 20201014

entity memory is
    port (
        
        );
end entity;

architecture behaviour of memory is


begin

end architecture;